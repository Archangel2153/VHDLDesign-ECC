-- include the STD_LOGIC_1164 package in the IEEE library for basic functionality
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- include the NUMERIC_STD package for arithmetic operations
use IEEE.NUMERIC_STD.ALL;

entity ecc_add_double is
    generic(
        n: integer := 8;
        log2n: integer := 3);
    port(
        start: in std_logic;
        rst: in std_logic;
        clk: in std_logic;
        add_double: in std_logic;
        busy: out std_logic;
        done: out std_logic;
        m_enable: in std_logic;
        m_din:in std_logic_vector(n-1 downto 0);
        m_dout:out std_logic_vector(n-1 downto 0);
        m_rw:in std_logic;
        m_address:in std_logic_vector(4 downto 0));
end ecc_add_double;

-- describe the behavior of the module in the architecture
architecture behavioral of ecc_add_double is

-- create the enumerated type 'my_state' to update and store the state of the FSM
type my_state is (s_idle, s_wait_ram, s_load_p, s_wait_p, s_load_add_1, s_add_1, s_write_add_1,
                  s_load_add_2, s_add_2, s_write_add_2,
						s_load_add_3, s_add_3, s_write_add_3,
						s_load_add_4, s_add_4, s_write_add_4,
						s_load_add_5, s_add_5, s_write_add_5,
						s_load_add_6, s_add_6, s_write_add_6,
						s_load_add_7, s_add_7, s_write_add_7,
						s_load_add_8, s_add_8, s_write_add_8,
						s_load_add_9, s_add_9, s_write_add_9,
						s_load_add_10, s_add_10, s_write_add_10,
						s_load_add_11, s_add_11, s_write_add_11,
						s_load_add_12, s_add_12, s_write_add_12,
						s_load_add_13, s_add_13, s_write_add_13,
						s_load_add_14, s_add_14, s_write_add_14,
						s_load_add_15, s_add_15, s_write_add_15,
						s_load_add_16, s_add_16, s_write_add_16,
						s_load_add_17, s_add_17, s_write_add_17,
						s_load_add_18, s_add_18, s_write_add_18,
						s_load_add_19, s_add_19, s_write_add_19,
						s_load_add_20, s_add_20, s_write_add_20,
						s_load_add_21, s_add_21, s_write_add_21,
						s_load_add_22, s_add_22, s_write_add_22,
						s_load_add_23, s_add_23, s_write_add_23,
						s_load_add_24, s_add_24, s_write_add_24,
						s_load_add_25, s_add_25, s_write_add_25,
						s_load_add_26, s_add_26, s_write_add_26,
						s_load_add_27, s_add_27, s_write_add_27,
						s_load_add_28, s_add_28, s_write_add_28,
						s_load_add_29, s_add_29, s_write_add_29,
						s_load_add_30, s_add_30, s_write_add_30,
						s_load_add_31, s_add_31, s_write_add_31,
						s_load_add_32, s_add_32, s_write_add_32,
						s_load_add_33, s_add_33, s_write_add_33,
						s_load_add_34, s_add_34, s_write_add_34,
						s_load_add_35, s_add_35, s_write_add_35,
						s_load_add_36, s_add_36, s_write_add_36,
						s_load_add_37, s_add_37, s_write_add_37,
						s_load_add_38, s_add_38, s_write_add_38,
						s_load_add_39, s_add_39, s_write_add_39,
						s_load_add_40, s_add_40, s_write_add_40,
						s_load_add_41, s_add_41, s_write_add_41,
						s_load_add_42, s_add_42, s_write_add_42,
						s_load_add_43, s_add_43, s_write_add_43,
						s_load_double_1, s_double_1, s_write_double_1,
						s_load_double_2, s_double_2, s_write_double_2,
						s_load_double_3, s_double_3, s_write_double_3,
						s_load_double_4, s_double_4, s_write_double_4,
						s_load_double_5, s_double_5, s_write_double_5,
						s_load_double_6, s_double_6, s_write_double_6,
						s_load_double_7, s_double_7, s_write_double_7,
						s_load_double_8, s_double_8, s_write_double_8,
						s_load_double_9, s_double_9, s_write_double_9,
						s_load_double_10, s_double_10, s_write_double_10,
						s_load_double_11, s_double_11, s_write_double_11,
						s_load_double_12, s_double_12, s_write_double_12,
						s_load_double_13, s_double_13, s_write_double_13,
						s_load_double_14, s_double_14, s_write_double_14,
						s_load_double_15, s_double_15, s_write_double_15,
						s_load_double_16, s_double_16, s_write_double_16,
						s_load_double_17, s_double_17, s_write_double_17,
						s_load_double_18, s_double_18, s_write_double_18,
						s_load_double_19, s_double_19, s_write_double_19,
						s_load_double_20, s_double_20, s_write_double_20,
						s_load_double_21, s_double_21, s_write_double_21,
						s_load_double_22, s_double_22, s_write_double_22,
						s_load_double_23, s_double_23, s_write_double_23,
						s_load_double_24, s_double_24, s_write_double_24,
						s_load_double_25, s_double_25, s_write_double_25,
						s_load_double_26, s_double_26, s_write_double_26,
						s_load_double_27, s_double_27, s_write_double_27,
						s_load_double_28, s_double_28, s_write_double_28,
						s_load_double_29, s_double_29, s_write_double_29,
						s_load_double_30, s_double_30, s_write_double_30,
						s_load_double_31, s_double_31, s_write_double_31,
						s_load_double_32, s_double_32, s_write_double_32,
						s_load_double_33, s_double_33, s_write_double_33,
						s_load_double_34, s_double_34, s_write_double_34,
						s_done);

-- declare internal signals
signal oper_o, oper_a, oper_b, address_i_1, address_i_2: std_logic_vector(4 downto 0);
signal a, b, p, product, din_i_1: std_logic_vector(n-1 downto 0);
signal state: my_state;
signal cmd: std_logic_vector(2 downto 0);
signal free, rw, enable, p_enable, a_start, a_done, rw_i, enable_i: std_logic;

-- declare the modarithn component
component modarithn
    generic(
        n: integer := 8;
		  log2n: integer := 3);
    port(
        a, b, p: in std_logic_vector(n-1 downto 0);
        rst, clk, start: in std_logic;
		  command: in std_logic_vector(1 downto 0);
        product: out std_logic_vector(n-1 downto 0);
        done: out std_logic);
end component;

-- declare the ram_double component
component ram_double
    generic(
        ws: integer := 8;
        ads: integer := 5);
    port(
        enable, clk, rw: in std_logic;
        din_a: in std_logic_vector((ws - 1) downto 0);
		  address_a, address_b: in std_logic_vector((ads - 1) downto 0);
        dout_a, dout_b: out std_logic_vector((ws - 1) downto 0));
end component;

begin

-- instantiate the modarithn component
-- map the generic parameter in the top design to the generic parameter in the component  
-- map the signals in the top design to the ports of the component
inst_modarithn: modarithn
    generic map(n => n,
	 log2n => log2n)
    port map(   a => a,
                b => b,
                p => p,
					 rst => rst,
					 clk => clk,
					 start => a_start,
					 command => cmd(1 downto 0),
                product => product,
                done => a_done);
					 
-- instantiate the ram_double component
-- map the generic parameter in the top design to the generic parameter in the component  
-- map the signals in the top design to the ports of the component
inst_ram_double: ram_double
    generic map(ws => n)
    port map(   enable => enable_i,
                clk => clk,
                rw => rw_i,
                din_a => din_i_1,
                address_a => address_i_2,
					 address_b => oper_b,
					 dout_a => a,
					 dout_b => b);

-- create the first multiplexer which selects between oper_a_address and oper_o_address					 
mux_1: process(oper_a, oper_o, rw)
begin
    if rw = '0' then
        address_i_1 <= oper_a;
    else
        address_i_1 <= oper_o;
    end if;
end process;

-- create the second multiplexer which selects between address_i_1 and m_address					 
mux_2: process(address_i_1, m_address, free)
begin
    if free = '0' then
        address_i_2 <= address_i_1;
    else
        address_i_2 <= m_address;
    end if;
end process;

-- create the third multiplexer which selects between m_din and product
mux_3: process(product, m_din, free)
begin
    if free = '0' then
        din_i_1 <= product;
    else
        din_i_1 <= m_din;
    end if;
end process;

-- create the fourth multiplexer which selects between rw and m_rw
mux_4: process(rw, m_rw, free)
begin
    if free = '0' then
        rw_i <= rw;
    else
        rw_i <= m_rw;
    end if;
end process;

-- create the fifth multiplexer which selects between enable and m_enable
mux_5: process(enable, m_enable, free)
begin
    if free = '0' then
        enable_i <= enable;
    else
        enable_i <= m_enable;
    end if;
end process;

-- store the value of 'b' in the register 'p' if 'p_enable' is '1' 
reg_p: process(clk)
begin
    if rising_edge(clk) then
        if p_enable = '1' then
            p <= b;
        end if;
    end if;
end process;

busy <= not(free);
m_dout <= a;

-- update and store the state of the FSM
-- (we lose 1 cycle by resetting the product register when the start signal comes)
FSM_state: process(rst, clk)
begin
    if rst = '1' then
        state <= s_idle;
    elsif rising_edge(clk) then
        case state is
            when s_idle =>
                if start = '1' then
                    state <= s_wait_ram;
                end if;
				when s_wait_ram =>
					 state <= s_load_p;
            when s_load_p =>
                state <= s_wait_p;
				when s_wait_p =>
                if add_double = '0' then
                    state <= s_load_add_1;
				    else
					     state <= s_load_double_1;
					 end if;
				when s_load_add_1 =>
                state <= s_add_1;
				when s_add_1 =>
				    if a_done = '1' then
                    state <= s_write_add_1;
					 end if;
				when s_write_add_1 =>
				    state <= s_load_add_2;
				when s_load_add_2 =>
                state <= s_add_2;
				when s_add_2 =>
				    if a_done = '1' then
                    state <= s_write_add_2;
					 end if;
				when s_write_add_2 =>
				    state <= s_load_add_3;
				when s_load_add_3 =>
                state <= s_add_3;
				when s_add_3 =>
				    if a_done = '1' then
                    state <= s_write_add_3;
					 end if;
				when s_write_add_3 =>
				    state <= s_load_add_4;
				when s_load_add_4 =>
                state <= s_add_4;
				when s_add_4 =>
				    if a_done = '1' then
                    state <= s_write_add_4;
					 end if;
				when s_write_add_4 =>
				    state <= s_load_add_5;
			   when s_load_add_5 =>
                state <= s_add_5;
				when s_add_5 =>
				    if a_done = '1' then
                    state <= s_write_add_5;
					 end if;
				when s_write_add_5 =>
				    state <= s_load_add_6;
				when s_load_add_6 =>
                state <= s_add_6;
				when s_add_6 =>
				    if a_done = '1' then
                    state <= s_write_add_6;
					 end if;
				when s_write_add_6 =>
				    state <= s_load_add_7;
				when s_load_add_7 =>
                state <= s_add_7;
				when s_add_7 =>
				    if a_done = '1' then
                    state <= s_write_add_7;
					 end if;
				when s_write_add_7 =>
				    state <= s_load_add_8;
				when s_load_add_8 =>
                state <= s_add_8;
				when s_add_8 =>
				    if a_done = '1' then
                    state <= s_write_add_8;
					 end if;
				when s_write_add_8 =>
				    state <= s_load_add_9;
				when s_load_add_9 =>
                state <= s_add_9;
				when s_add_9 =>
				    if a_done = '1' then
                    state <= s_write_add_9;
					 end if;
				when s_write_add_9 =>
				    state <= s_load_add_10;
				when s_load_add_10 =>
                state <= s_add_10;
				when s_add_10 =>
				    if a_done = '1' then
                    state <= s_write_add_10;
					 end if;
				when s_write_add_10 =>
				    state <= s_load_add_11;
				when s_load_add_11 =>
                state <= s_add_11;
				when s_add_11 =>
				    if a_done = '1' then
                    state <= s_write_add_11;
					 end if;
				when s_write_add_11 =>
				    state <= s_load_add_12;
				when s_load_add_12 =>
                state <= s_add_12;
				when s_add_12 =>
				    if a_done = '1' then
                    state <= s_write_add_12;
					 end if;
				when s_write_add_12 =>
				    state <= s_load_add_13;
				when s_load_add_13 =>
                state <= s_add_13;
				when s_add_13 =>
				    if a_done = '1' then
                    state <= s_write_add_13;
					 end if;
				when s_write_add_13 =>
				    state <= s_load_add_14;
				when s_load_add_14 =>
                state <= s_add_14;
				when s_add_14 =>
				    if a_done = '1' then
                    state <= s_write_add_14;
					 end if;
				when s_write_add_14 =>
				    state <= s_load_add_15;
				when s_load_add_15 =>
                state <= s_add_15;
				when s_add_15 =>
				    if a_done = '1' then
                    state <= s_write_add_15;
					 end if;
				when s_write_add_15 =>
				    state <= s_load_add_16;
				when s_load_add_16 =>
                state <= s_add_16;
				when s_add_16 =>
				    if a_done = '1' then
                    state <= s_write_add_16;
					 end if;
				when s_write_add_16 =>
				    state <= s_load_add_17;
				when s_load_add_17 =>
                state <= s_add_17;
				when s_add_17 =>
				    if a_done = '1' then
                    state <= s_write_add_17;
					 end if;
				when s_write_add_17 =>
				    state <= s_load_add_18;
				when s_load_add_18 =>
                state <= s_add_18;
				when s_add_18 =>
				    if a_done = '1' then
                    state <= s_write_add_18;
					 end if;
				when s_write_add_18 =>
				    state <= s_load_add_19;
				when s_load_add_19 =>
                state <= s_add_19;
				when s_add_19 =>
				    if a_done = '1' then
                    state <= s_write_add_19;
					 end if;
				when s_write_add_19 =>
				    state <= s_load_add_20;
				when s_load_add_20 =>
                state <= s_add_20;
				when s_add_20 =>
				    if a_done = '1' then
                    state <= s_write_add_20;
					 end if;
				when s_write_add_20 =>
				    state <= s_load_add_21;
				when s_load_add_21 =>
                state <= s_add_21;
				when s_add_21 =>
				    if a_done = '1' then
                    state <= s_write_add_21;
					 end if;
				when s_write_add_21 =>
				    state <= s_load_add_22;
				when s_load_add_22 =>
                state <= s_add_22;
				when s_add_22 =>
				    if a_done = '1' then
                    state <= s_write_add_22;
					 end if;
				when s_write_add_22 =>
				    state <= s_load_add_23;
				when s_load_add_23 =>
                state <= s_add_23;
				when s_add_23 =>
				    if a_done = '1' then
                    state <= s_write_add_23;
					 end if;
				when s_write_add_23 =>
				    state <= s_load_add_24;
				when s_load_add_24 =>
                state <= s_add_24;
				when s_add_24 =>
				    if a_done = '1' then
                    state <= s_write_add_24;
					 end if;
				when s_write_add_24 =>
				    state <= s_load_add_25;
				when s_load_add_25 =>
                state <= s_add_25;
				when s_add_25 =>
				    if a_done = '1' then
                    state <= s_write_add_25;
					 end if;
				when s_write_add_25 =>
				    state <= s_load_add_26;
				when s_load_add_26 =>
                state <= s_add_26;
				when s_add_26 =>
				    if a_done = '1' then
                    state <= s_write_add_26;
					 end if;
				when s_write_add_26 =>
				    state <= s_load_add_27;
				when s_load_add_27 =>
                state <= s_add_27;
				when s_add_27 =>
				    if a_done = '1' then
                    state <= s_write_add_27;
					 end if;
				when s_write_add_27 =>
				    state <= s_load_add_28;
				when s_load_add_28 =>
                state <= s_add_28;
				when s_add_28 =>
				    if a_done = '1' then
                    state <= s_write_add_28;
					 end if;
				when s_write_add_28 =>
				    state <= s_load_add_29;
				when s_load_add_29 =>
                state <= s_add_29;
				when s_add_29 =>
				    if a_done = '1' then
                    state <= s_write_add_29;
					 end if;
				when s_write_add_29 =>
				    state <= s_load_add_30;
				when s_load_add_30 =>
                state <= s_add_30;
				when s_add_30 =>
				    if a_done = '1' then
                    state <= s_write_add_30;
					 end if;
				when s_write_add_30 =>
				    state <= s_load_add_31;
				when s_load_add_31 =>
                state <= s_add_31;
				when s_add_31 =>
				    if a_done = '1' then
                    state <= s_write_add_31;
					 end if;
				when s_write_add_31 =>
				    state <= s_load_add_32;
				when s_load_add_32 =>
                state <= s_add_32;
				when s_add_32 =>
				    if a_done = '1' then
                    state <= s_write_add_32;
					 end if;
				when s_write_add_32 =>
				    state <= s_load_add_33;
			   when s_load_add_33 =>
                state <= s_add_33;
				when s_add_33 =>
				    if a_done = '1' then
                    state <= s_write_add_33;
					 end if;
				when s_write_add_33 =>
				    state <= s_load_add_34;
			   when s_load_add_34 =>
                state <= s_add_34;
				when s_add_34 =>
				    if a_done = '1' then
                    state <= s_write_add_34;
					 end if;
				when s_write_add_34 =>
				    state <= s_load_add_35;
				when s_load_add_35 =>
                state <= s_add_35;
				when s_add_35 =>
				    if a_done = '1' then
                    state <= s_write_add_35;
					 end if;
				when s_write_add_35 =>
				    state <= s_load_add_36;
				when s_load_add_36 =>
                state <= s_add_36;
				when s_add_36 =>
				    if a_done = '1' then
                    state <= s_write_add_36;
					 end if;
				when s_write_add_36 =>
				    state <= s_load_add_37;
				when s_load_add_37 =>
                state <= s_add_37;
				when s_add_37 =>
				    if a_done = '1' then
                    state <= s_write_add_37;
					 end if;
				when s_write_add_37 =>
				    state <= s_load_add_38;
				when s_load_add_38 =>
                state <= s_add_38;
				when s_add_38 =>
				    if a_done = '1' then
                    state <= s_write_add_38;
					 end if;
				when s_write_add_38 =>
				    state <= s_load_add_39;
				when s_load_add_39 =>
                state <= s_add_39;
				when s_add_39 =>
				    if a_done = '1' then
                    state <= s_write_add_39;
					 end if;
				when s_write_add_39 =>
				    state <= s_load_add_40;
				when s_load_add_40 =>
                state <= s_add_40;
				when s_add_40 =>
				    if a_done = '1' then
                    state <= s_write_add_40;
					 end if;
				when s_write_add_40 =>
				    state <= s_load_add_41;
				when s_load_add_41 =>
                state <= s_add_41;
				when s_add_41 =>
				    if a_done = '1' then
                    state <= s_write_add_41;
					 end if;
				when s_write_add_41 =>
				    state <= s_load_add_42;
				when s_load_add_42 =>
                state <= s_add_42;
				when s_add_42 =>
				    if a_done = '1' then
                    state <= s_write_add_42;
					 end if;
				when s_write_add_42 =>
				    state <= s_load_add_43;
				when s_load_add_43 =>
                state <= s_add_43;
				when s_add_43 =>
				    if a_done = '1' then
                    state <= s_write_add_43;
					 end if;
				when s_write_add_43 =>
				    state <= s_done;
				when s_load_double_1 =>
                state <= s_double_1;
				when s_double_1 =>
				    if a_done = '1' then
                    state <= s_write_double_1;
					 end if;
				when s_write_double_1 =>
				    state <= s_load_double_2;
				when s_load_double_2 =>
                state <= s_double_2;
				when s_double_2 =>
				    if a_done = '1' then
                    state <= s_write_double_2;
					 end if;
				when s_write_double_2 =>
				    state <= s_load_double_3;
				when s_load_double_3 =>
                state <= s_double_3;
				when s_double_3 =>
				    if a_done = '1' then
                    state <= s_write_double_3;
					 end if;
				when s_write_double_3 =>
				    state <= s_load_double_4;
				when s_load_double_4 =>
                state <= s_double_4;
				when s_double_4 =>
				    if a_done = '1' then
                    state <= s_write_double_4;
					 end if;
				when s_write_double_4 =>
				    state <= s_load_double_5;
			   when s_load_double_5 =>
                state <= s_double_5;
				when s_double_5 =>
				    if a_done = '1' then
                    state <= s_write_double_5;
					 end if;
				when s_write_double_5 =>
				    state <= s_load_double_6;
				when s_load_double_6 =>
                state <= s_double_6;
				when s_double_6 =>
				    if a_done = '1' then
                    state <= s_write_double_6;
					 end if;
				when s_write_double_6 =>
				    state <= s_load_double_7;
				when s_load_double_7 =>
                state <= s_double_7;
				when s_double_7 =>
				    if a_done = '1' then
                    state <= s_write_double_7;
					 end if;
				when s_write_double_7 =>
				    state <= s_load_double_8;
				when s_load_double_8 =>
                state <= s_double_8;
				when s_double_8 =>
				    if a_done = '1' then
                    state <= s_write_double_8;
					 end if;
				when s_write_double_8 =>
				    state <= s_load_double_9;
				when s_load_double_9 =>
                state <= s_double_9;
				when s_double_9 =>
				    if a_done = '1' then
                    state <= s_write_double_9;
					 end if;
				when s_write_double_9 =>
				    state <= s_load_double_10;
				when s_load_double_10 =>
                state <= s_double_10;
				when s_double_10 =>
				    if a_done = '1' then
                    state <= s_write_double_10;
					 end if;
				when s_write_double_10 =>
				    state <= s_load_double_11;
				when s_load_double_11 =>
                state <= s_double_11;
				when s_double_11 =>
				    if a_done = '1' then
                    state <= s_write_double_11;
					 end if;
				when s_write_double_11 =>
				    state <= s_load_double_12;
				when s_load_double_12 =>
                state <= s_double_12;
				when s_double_12 =>
				    if a_done = '1' then
                    state <= s_write_double_12;
					 end if;
				when s_write_double_12 =>
				    state <= s_load_double_13;
				when s_load_double_13 =>
                state <= s_double_13;
				when s_double_13 =>
				    if a_done = '1' then
                    state <= s_write_double_13;
					 end if;
				when s_write_double_13 =>
				    state <= s_load_double_14;
				when s_load_double_14 =>
                state <= s_double_14;
				when s_double_14 =>
				    if a_done = '1' then
                    state <= s_write_double_14;
					 end if;
				when s_write_double_14 =>
				    state <= s_load_double_15;
				when s_load_double_15 =>
                state <= s_double_15;
				when s_double_15 =>
				    if a_done = '1' then
                    state <= s_write_double_15;
					 end if;
				when s_write_double_15 =>
				    state <= s_load_double_16;
				when s_load_double_16 =>
                state <= s_double_16;
				when s_double_16 =>
				    if a_done = '1' then
                    state <= s_write_double_16;
					 end if;
				when s_write_double_16 =>
				    state <= s_load_double_17;
				when s_load_double_17 =>
                state <= s_double_17;
				when s_double_17 =>
				    if a_done = '1' then
                    state <= s_write_double_17;
					 end if;
				when s_write_double_17 =>
				    state <= s_load_double_18;
				when s_load_double_18 =>
                state <= s_double_18;
				when s_double_18 =>
				    if a_done = '1' then
                    state <= s_write_double_18;
					 end if;
				when s_write_double_18 =>
				    state <= s_load_double_19;
				when s_load_double_19 =>
                state <= s_double_19;
				when s_double_19 =>
				    if a_done = '1' then
                    state <= s_write_double_19;
					 end if;
				when s_write_double_19 =>
				    state <= s_load_double_20;
				when s_load_double_20 =>
                state <= s_double_20;
				when s_double_20 =>
				    if a_done = '1' then
                    state <= s_write_double_20;
					 end if;
				when s_write_double_20 =>
				    state <= s_load_double_21;
				when s_load_double_21 =>
                state <= s_double_21;
				when s_double_21 =>
				    if a_done = '1' then
                    state <= s_write_double_21;
					 end if;
				when s_write_double_21 =>
				    state <= s_load_double_22;
				when s_load_double_22 =>
                state <= s_double_22;
				when s_double_22 =>
				    if a_done = '1' then
                    state <= s_write_double_22;
					 end if;
				when s_write_double_22 =>
				    state <= s_load_double_23;
				when s_load_double_23 =>
                state <= s_double_23;
				when s_double_23 =>
				    if a_done = '1' then
                    state <= s_write_double_23;
					 end if;
				when s_write_double_23 =>
				    state <= s_load_double_24;
				when s_load_double_24 =>
                state <= s_double_24;
				when s_double_24 =>
				    if a_done = '1' then
                    state <= s_write_double_24;
					 end if;
				when s_write_double_24 =>
				    state <= s_load_double_25;
				when s_load_double_25 =>
                state <= s_double_25;
				when s_double_25 =>
				    if a_done = '1' then
                    state <= s_write_double_25;
					 end if;
				when s_write_double_25 =>
				    state <= s_load_double_26;
				when s_load_double_26 =>
                state <= s_double_26;
				when s_double_26 =>
				    if a_done = '1' then
                    state <= s_write_double_26;
					 end if;
				when s_write_double_26 =>
				    state <= s_load_double_27;
				when s_load_double_27 =>
                state <= s_double_27;
				when s_double_27 =>
				    if a_done = '1' then
                    state <= s_write_double_27;
					 end if;
				when s_write_double_27 =>
				    state <= s_load_double_28;
				when s_load_double_28 =>
                state <= s_double_28;
				when s_double_28 =>
				    if a_done = '1' then
                    state <= s_write_double_28;
					 end if;
				when s_write_double_28 =>
				    state <= s_load_double_29;
				when s_load_double_29 =>
                state <= s_double_29;
				when s_double_29 =>
				    if a_done = '1' then
                    state <= s_write_double_29;
					 end if;
				when s_write_double_29 =>
				    state <= s_load_double_30;
				when s_load_double_30 =>
                state <= s_double_30;
				when s_double_30 =>
				    if a_done = '1' then
                    state <= s_write_double_30;
					 end if;
				when s_write_double_30 =>
				    state <= s_load_double_31;
				when s_load_double_31 =>
                state <= s_double_31;
				when s_double_31 =>
				    if a_done = '1' then
                    state <= s_write_double_31;
					 end if;
				when s_write_double_31 =>
				    state <= s_load_double_32;
				when s_load_double_32 =>
                state <= s_double_32;
				when s_double_32 =>
				    if a_done = '1' then
                    state <= s_write_double_32;
					 end if;
				when s_write_double_32 =>
				    state <= s_load_double_33;
			   when s_load_double_33 =>
                state <= s_double_33;
				when s_double_33 =>
				    if a_done = '1' then
                    state <= s_write_double_33;
					 end if;
				when s_write_double_33 =>
				    state <= s_load_double_34;
			   when s_load_double_34 =>
                state <= s_double_34;
				when s_double_34 =>
				    if a_done = '1' then
                    state <= s_write_double_34;
					 end if;
				when s_write_double_34 =>
				    state <= s_done;
            when others =>
                state <= s_idle;
        end case;
    end if;
end process;

FSM_out: process(state)
begin
    case state is
        when s_idle =>
		      oper_a <= std_logic_vector(to_unsigned(31, 5));
				oper_b <= std_logic_vector(to_unsigned(31, 5));
				oper_o <= std_logic_vector(to_unsigned(31, 5));
				cmd <= std_logic_vector(to_unsigned(7, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '1';
		  when s_wait_ram =>
            oper_a <= std_logic_vector(to_unsigned(31, 5));
				oper_b <= std_logic_vector(to_unsigned(0, 5));
				oper_o <= std_logic_vector(to_unsigned(31, 5));
				cmd <= std_logic_vector(to_unsigned(7, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when s_load_p =>
		      oper_a <= std_logic_vector(to_unsigned(31, 5));
				oper_b <= std_logic_vector(to_unsigned(0, 5));
				oper_o <= std_logic_vector(to_unsigned(31, 5));
				cmd <= std_logic_vector(to_unsigned(6, 3));
				p_enable <= '1';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_wait_p =>
		      oper_a <= std_logic_vector(to_unsigned(31, 5));
				oper_b <= std_logic_vector(to_unsigned(31, 5));
				oper_o <= std_logic_vector(to_unsigned(31, 5));
				cmd <= std_logic_vector(to_unsigned(7, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_load_add_1 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(6, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_1 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(6, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_1 =>
				oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(6, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_2 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(7, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_2 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(7, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_2 =>
				oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(7, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_3 =>
		      oper_a <= std_logic_vector(to_unsigned(5, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_3 =>
		      oper_a <= std_logic_vector(to_unsigned(5, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_3 =>
				oper_a <= std_logic_vector(to_unsigned(5, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_4 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_4 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_4 =>
				oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_5 =>
		      oper_a <= std_logic_vector(to_unsigned(6, 5));
				oper_b <= std_logic_vector(to_unsigned(7, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_5 =>
		      oper_a <= std_logic_vector(to_unsigned(6, 5));
				oper_b <= std_logic_vector(to_unsigned(7, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_5 =>
				oper_a <= std_logic_vector(to_unsigned(6, 5));
				oper_b <= std_logic_vector(to_unsigned(7, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_6 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(16, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_6 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(16, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_6 =>
				oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(16, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_7 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_7 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_7 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_8 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(16, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_8 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(16, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_8 =>
				oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(16, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_9 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_9 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_9 =>
				oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_10 =>
		      oper_a <= std_logic_vector(to_unsigned(7, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_10 =>
		      oper_a <= std_logic_vector(to_unsigned(7, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_10 =>
				oper_a <= std_logic_vector(to_unsigned(7, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_11 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_11 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_11 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_12 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_12 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_12 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_13 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_13 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_13 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_14 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_14 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_14 =>
				oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_15 =>
		      oper_a <= std_logic_vector(to_unsigned(6, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_15 =>
		      oper_a <= std_logic_vector(to_unsigned(6, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_15 =>
				oper_a <= std_logic_vector(to_unsigned(6, 5));
				oper_b <= std_logic_vector(to_unsigned(8, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_16 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_16 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_16 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_17 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_17 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_17 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_18 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_18 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_18 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';	
			when s_load_add_19 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_19 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_19 =>
				oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
			when s_load_add_20 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_20 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_20 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when s_load_add_21 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_21 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_21 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_22 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_22 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_22 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when s_load_add_23 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_23 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_23 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when s_load_add_24 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_24 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_24 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when s_load_add_25 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_25 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_25 =>
				oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when s_load_add_26 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_26 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_26 =>
				oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_27 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_27 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_27 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_28 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_28 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_28 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_29 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_29 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_29 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_30 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_30 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_30 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_31 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_31 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_31 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_32 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_32 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_32 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_33 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_33 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_33 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_34 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_34 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_34 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_35 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_35 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_35 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_36 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_36 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_36 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_37 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_37 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_37 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_38 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(10, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_38 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(10, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_38 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(10, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_39 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_39 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_39 =>
				oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_40 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(9, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_40 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(9, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_40 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(9, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_41 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_41 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_41 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(19, 5));
				oper_o <= std_logic_vector(to_unsigned(19, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_42 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_42 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_42 =>
				oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_add_43 =>
		      oper_a <= std_logic_vector(to_unsigned(19, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(11, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_add_43 =>
		      oper_a <= std_logic_vector(to_unsigned(19, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(11, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_add_43 =>
				oper_a <= std_logic_vector(to_unsigned(19, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(11, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_1 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(3, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_1 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(3, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_1 =>
				oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(3, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_2 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_2 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_2 =>
				oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(13, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_3 =>
		      oper_a <= std_logic_vector(to_unsigned(5, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_3 =>
		      oper_a <= std_logic_vector(to_unsigned(5, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_3 =>
				oper_a <= std_logic_vector(to_unsigned(5, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_4 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_4 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_4 =>
				oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(4, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_5 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_5 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_5 =>
				oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_6 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_6 =>
		      oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_6 =>
				oper_a <= std_logic_vector(to_unsigned(3, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_7 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_7 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_7 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_8 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_8 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_8 =>
				oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_9 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_9 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_9 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_10 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_10 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_10 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_11 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_11 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_11 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_12 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_12 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_12 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_13 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_13 =>
		      oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_13 =>
				oper_a <= std_logic_vector(to_unsigned(13, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_14 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_14 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_14 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(17, 5));
				oper_o <= std_logic_vector(to_unsigned(17, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_15 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_15 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_15 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(16, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_16 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_16 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_16 =>
				oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_17 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_17 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_17 =>
				oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_18 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_18 =>
		      oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_18 =>
				oper_a <= std_logic_vector(to_unsigned(2, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_19 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_19 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_19 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_20 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_20 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_20 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_21 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_21 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_21 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_22 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_22 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_22 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(15, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_23 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_23 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_23 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(15, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_24 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_24 =>
		      oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_24 =>
				oper_a <= std_logic_vector(to_unsigned(15, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_25 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_25 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_25 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_26 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_26 =>
		      oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_26 =>
				oper_a <= std_logic_vector(to_unsigned(12, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(12, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_27 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_27 =>
		      oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_27 =>
				oper_a <= std_logic_vector(to_unsigned(4, 5));
				oper_b <= std_logic_vector(to_unsigned(5, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_28 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_28 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_28 =>
				oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(14, 5));
				oper_o <= std_logic_vector(to_unsigned(14, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_29 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(10, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_29 =>
		      oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(10, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_29 =>
				oper_a <= std_logic_vector(to_unsigned(17, 5));
				oper_b <= std_logic_vector(to_unsigned(12, 5));
				oper_o <= std_logic_vector(to_unsigned(10, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_30 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_30 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_30 =>
				oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_31 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(9, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_31 =>
		      oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(9, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_31 =>
				oper_a <= std_logic_vector(to_unsigned(16, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(9, 5));
				cmd <= std_logic_vector(to_unsigned(1, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_32 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_32 =>
		      oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_32 =>
				oper_a <= std_logic_vector(to_unsigned(14, 5));
				oper_b <= std_logic_vector(to_unsigned(13, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(3, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_33 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_33 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_33 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(18, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
		  when s_load_double_34 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(11, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '1';
				enable <= '1';
		      free <= '0';
		  when s_double_34 =>
		      oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(11, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '0';
				a_start <= '0';
				enable <= '0';
		      free <= '0';
		  when s_write_double_34 =>
				oper_a <= std_logic_vector(to_unsigned(18, 5));
				oper_b <= std_logic_vector(to_unsigned(18, 5));
				oper_o <= std_logic_vector(to_unsigned(11, 5));
				cmd <= std_logic_vector(to_unsigned(0, 3));
				p_enable <= '0';
				done <= '0';
				rw <= '1';
				a_start <= '0';
				enable <= '1';
		      free <= '0';
        when others =>
		      oper_a <= std_logic_vector(to_unsigned(31, 5));
				oper_b <= std_logic_vector(to_unsigned(31, 5));
				oper_o <= std_logic_vector(to_unsigned(31, 5));
				cmd <= std_logic_vector(to_unsigned(7, 3));
            free <= '0';
				done <= '1';
				rw <= '0';
            enable <= '0';
				a_start <= '0';
				p_enable <= '0';
    end case;
end process;

end behavioral;
